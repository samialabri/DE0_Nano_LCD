library verilog;
use verilog.vl_types.all;
entity teshBench is
end teshBench;
